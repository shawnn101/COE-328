library verilog;
use verilog.vl_types.all;
entity CombinedASU1_vlg_vec_tst is
end CombinedASU1_vlg_vec_tst;
