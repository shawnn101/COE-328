library verilog;
use verilog.vl_types.all;
entity decodeModified_vlg_vec_tst is
end decodeModified_vlg_vec_tst;
