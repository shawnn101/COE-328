library verilog;
use verilog.vl_types.all;
entity ASU_vlg_vec_tst is
end ASU_vlg_vec_tst;
