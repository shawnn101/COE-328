library verilog;
use verilog.vl_types.all;
entity CombinedASU2_vlg_vec_tst is
end CombinedASU2_vlg_vec_tst;
