library verilog;
use verilog.vl_types.all;
entity sseg_vlg_vec_tst is
end sseg_vlg_vec_tst;
